// Things to test :

// - Read / Write (normal)
// - Test TREADY and TVILID outputs when full and empty
// - Test R/W when both S & M want infos
// - Test TLAST handling